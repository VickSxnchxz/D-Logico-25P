entity p1 is 
port(
	a: in bit;
	c: out bit
);
end p1;

architecture arch_p1 of p1 is
	begin 
		c <= a;
end arch_p1;
		